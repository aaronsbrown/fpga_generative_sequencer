package proj_defs_pkg;

    // Define parameters, types, enums, structs here
    // Example:
    // parameter DATA_WIDTH = 8;
    // typedef logic [DATA_WIDTH-1:0] data_t;

endpackage : proj_defs_pkg